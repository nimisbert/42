* Circuit :
* Photovoltaic Cell Model
.model pvcell D (
+ Is=10n
+ Rs=.5
+ N=77.06
+ Cjo=10n
+ M=.5
+ Eg=85
+ Xti=230
+ BV=30
+ IBV=.001
+ Vj=.4
+ Iave=1
+ Vpk=30
+ mfg=Generic
+ type=PV
+ )

.subckt pvpanel A K
I1 K A {Il}
D1 A K pvcell Is={Is} Imax={Im} Vmax={Vm} N={Vm}*38.6/log({Im}/{Is}) XTI=3*{N} EG=1.11*{N}
.ends